library ieee;
use ieee.std_logic_1164.all;

entity mux4t1_N is
  generic (
    N : integer := 32  -- Width of the data inputs/outputs
  );
  port (
    i_sel  : in  std_logic_vector(1 downto 0); -- 2-bit select
    i_D0   : in  std_logic_vector(N-1 downto 0);
    i_D1   : in  std_logic_vector(N-1 downto 0);
    i_D2   : in  std_logic_vector(N-1 downto 0);
    i_D3   : in  std_logic_vector(N-1 downto 0);
    o_O    : out std_logic_vector(N-1 downto 0)
  );
end mux4t1_N;

architecture Behavioral of mux4t1_N is
begin
  -- Select signal based on i_sel
  process(i_sel, i_D0, i_D1, i_D2, i_D3)
  begin
    case i_sel is
      when "00" => o_O <= i_D0;
      when "01" => o_O <= i_D1;
      when "10" => o_O <= i_D2;
      when "11" => o_O <= i_D3;
      when others => o_O <= (others => '0'); -- If no option selected, default is 0x0
    end case;
  end process;
end Behavioral;
